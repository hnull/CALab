module Data_memory(input [31:0]address,write_data,input mem_read,mem_write,input clk,rst,output [31:0] read_data);
  reg [31:0] memory [6500:0];
  assign read_data = mem_read ? memory[address] : 32'b0;

  always @ ( posedge clk ) begin
    if (mem_write) begin
      memory[address] = write_data;
    end
     // memory[1000] = 32'b00000000000000000000000000000001;
     // memory[1004] = 32'b00000000000000000000000000000010;
     // memory[1008] = 32'b00000000000000000000000000000011;
     // memory[1012] = 32'b00000000000000000000000000000100;
     // memory[1016] = 32'b00000000000000000000000000000101;
     // memory[1020] = 32'b00000000000000000000000000000110;
     // memory[1024] = 32'b00000000000000000000000000000111;
     // memory[1028] = 32'b00000000000000000000000000001000;
     // memory[1032] = 32'b00000000000000000000000000001001;
     // memory[1036] = 32'b00000000000000000000000000001010;
     // memory[1040] = 32'b00000000000000000000000000001011;
     // memory[1044] = 32'b00000000000000000000000000001100;
     // memory[1048] = 32'b00000000000000000000000000001101;
     // memory[1052] = 32'b00000000000000000000000000001110;
     // memory[1056] = 32'b00000000000000000000000000001111;
     // memory[1060] = 32'b00000000000000000000000000010000;
     // memory[1064] = 32'b00000000000000000000000000010001;
     // memory[1068] = 32'b00000000000000000000000000010010;
     // memory[1072] = 32'b00000000000000000000000000010011;
     // memory[1076] = 32'b00000000000000000000000000010100;
  end

endmodule //data_memory
