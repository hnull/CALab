module Instruction
  (
    input[31:0] adrs,
    output[31:0] inst
  );

  wire [31:0] Mem [100:0];

  assign Mem[0] = 32'b00000000000000000000000000000000;
  assign Mem[4] = 32'b10000000000000010000011000001010;
  assign Mem[8] = 32'b00000100000000010001000000000000;
  assign Mem[12] = 32'b00001100000000010001100000000000;
  assign Mem[16] = 32'b00010100010000110010000000000000;
  assign Mem[20] = 32'b10000100011001010001101000110100;
  assign Mem[24] = 32'b00011000011001000010100000000000;
  assign inst = Mem[adrs];

endmodule
